//
// The Test Bench File for 
// Thunderbird Turn Signal
// 
// Neil Nie
// (c) 2018, All Rights Reserved
//


module tb ();

//	logic clk, reset;
//	logic left, right;
//	logic LA, LB, LC, RA, RB, RC;

endmodule
